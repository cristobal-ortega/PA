LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FETCH IS 
	PORT (clock : IN	STD_LOGIC;
			inst  : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000");

END FETCH;


ARCHITECTURE Structure OF FETCH IS
BEGIN

END Structure;