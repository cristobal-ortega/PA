amspodnaspdnaspd