LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY EXECUTION1 IS 
	PORT (clock : IN	STD_LOGIC;
			op  : IN STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
			w	 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000");

END EXECUTION1;


ARCHITECTURE Structure OF EXECUTION1 IS
BEGIN

END Structure;