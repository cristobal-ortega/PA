LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

ENTITY suchControl IS 
	PORT (clock : IN	STD_LOGIC;

			);

END suchControl;


ARCHITECTURE Structure OF suchControl IS

--structural hazards
--data hazards
	
BEGIN

	PROCESS(clock)
	BEGIN

	END PROCESS;

END Structure;