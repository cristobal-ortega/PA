LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY MEMORY1_WRITEBACK IS 
	PORT (clock : IN	STD_LOGIC;
			data_in  : IN STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000";
			data_out	 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000");

END MEMORY1_WRITEBACK;


ARCHITECTURE Structure OF MEMORY1_WRITEBACK IS
BEGIN

END Structure;