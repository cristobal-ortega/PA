LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FETCH IS 
	PORT (clock : IN	STD_LOGIC);

END FETCH;


ARCHITECTURE Structure OF FETCH IS
BEGIN

END Structure;