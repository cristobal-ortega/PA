LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY DECODE1_EXECUTION1 IS 
	PORT (clock : IN	STD_LOGIC;
			op_in  : IN STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
			op_out : OUT STD_LOGIC_VECTOR(3 DOWNTO 0) :="0000");

END DECODE1_EXECUTION1;


ARCHITECTURE Structure OF DECODE1_EXECUTION1 IS
BEGIN

END Structure;