LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY MEMORY1 IS 
	PORT (clock : IN	STD_LOGIC;
	
			instr_in : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			op_in : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			w 		 : IN STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000";
			
			data	 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000";
			request	 : OUT STD_LOGIC := '0'
			);

END MEMORY1;


ARCHITECTURE Structure OF MEMORY1 IS
BEGIN

	data <= w;
END Structure;