LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY WRITEBACK IS 
	PORT (clock : IN	STD_LOGIC;
			data	: IN STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000";
			regwrite : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000");

END WRITEBACK;


ARCHITECTURE Structure OF WRITEBACK IS
BEGIN
	regwrite <= data;
END Structure;