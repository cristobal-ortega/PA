LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY D1 IS 
	PORT (clock : IN	STD_LOGIC);

END D1;


ARCHITECTURE Structure OF D1 IS
BEGIN

END Structure;