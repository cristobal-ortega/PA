LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FETCH_DECODE1 IS 
	PORT (clock : IN	STD_LOGIC);

END FETCH_DECODE1;


ARCHITECTURE Structure OF FETCH_DECODE1 IS
BEGIN

END Structure;