LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY DECODE1 IS 
	PORT (clock : IN	STD_LOGIC);

END DECODE1;


ARCHITECTURE Structure OF DECODE1 IS
BEGIN

END Structure;