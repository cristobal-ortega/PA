LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FETCH_D1 IS 
	PORT (clock : IN	STD_LOGIC);

END FETCH_D1;


ARCHITECTURE Structure OF FETCH_D1 IS
BEGIN

END Structure;