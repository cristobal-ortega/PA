LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY EXECUTION1_MEMORY1 IS 
	PORT (clock : IN	STD_LOGIC;
			w_in  : IN STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000";
			w_out	 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000");

END EXECUTION1_MEMORY1;


ARCHITECTURE Structure OF EXECUTION1_MEMORY1 IS
BEGIN

END Structure;