LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FETCH_DECODE1 IS 
	PORT (clock : IN	STD_LOGIC;
			inst_in  : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			inst_out : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000" );

END FETCH_DECODE1;


ARCHITECTURE Structure OF FETCH_DECODE1 IS
BEGIN

END Structure;